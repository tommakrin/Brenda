----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:47:48 04/27/2016 
-- Design Name: 
-- Module Name:    COMPARE_Unit - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.ALL;

entity COMPARE_Unit is

	port( POSITION	: in std_logic_vector(10 downto 0);
			SAD		: in std_logic_vector(15 downto 0);
			LOAD_EN	: in std_logic;
			CLK		: in std_logic;
			RESET		: in std_logic;
			MINPOS	: out std_logic_vector(10 downto 0)
			);

end COMPARE_Unit;

architecture Behavioral of COMPARE_Unit is

--Component Declaration
component X16Comparator is
	port (  
	  sad_cur, sad	: in std_logic_vector(15 downto 0);
	  pos_cur, pos	: in std_logic_vector(10 downto 0);
	  minSAD			: out std_logic_vector(15 downto 0);
	  minPOS			: out std_logic_vector(10 downto 0);
	  clk, rst : in std_logic
   );
end component;

component reg54 is
	generic (regCount : integer := 54);
	port ( clk : in std_logic;
			 rst : in std_logic;
			 loadEn : in std_logic;
			 reg_in : in std_logic_vector (regCount-1 downto 0);
			 reg_out : out std_logic_vector (regCount-1 downto 0)
			 );
end component;

signal reg_input:  std_logic_vector(53 downto 0);
signal reg_output: std_logic_vector(53 downto 0);
signal minPOS_int: std_logic_vector(10 downto 0);
signal minSAD_int: std_logic_vector(15 downto 0):= (others => '1');


begin
	minPOS <= minPOS_int;
	reg_input <= POSITION & SAD & minPOS_int & minSAD_int;
	
	COMP: X16Comparator port map(reg_output(42 downto 27), reg_output(15 downto 0),
										  reg_output(53 downto 43), reg_output(26 downto 16),
										  minSAD_int, minPOS_int, CLK, RESET);
	REG: reg54 port map(CLK, RESET, LOAD_EN, reg_input, reg_output);
	
end Behavioral;


